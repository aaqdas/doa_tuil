module basic_test(
    input   [7:0] i_a,
    input   [7:0] i_b,
    output  [7:0] o_c
);

assign o_c = i_a + i_b;

endmodule 